class AHB_master_monitor1 extends uvm_monitor;

endclass