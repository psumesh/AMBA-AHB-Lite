class AHB_monitor1 extends uvm_monitor;

endclass